//==============================================================================
// AU_incdec.v
//
// Incrementer-decrementer using parallel-prefix propagate-lookahead logic.
//------------------------------------------------------------------------------
// Copyright (c) 2023 Guangxi Liu
//
// This source code is licensed under the MIT license found in the
// LICENSE file in the root directory of this source tree.
//==============================================================================


module AU_incdec #(
    parameter integer WIDTH = 8,  // word length of input (>= 1)
    parameter integer ARCH  = 0   // architecture (0 to 2)
) (
    // Data interface
    input  [WIDTH-1:0] a,        // input data
    input              inc_dec,  // control, 0:increment, 1:decrement
    output [WIDTH-1:0] z         // increment or decrement
);


    // Structural model
    generate
        wire [WIDTH-1:0] at;
        wire [WIDTH-1:0] po;

        if (WIDTH == 1) begin : g_z_1
            // Calculate result bit
            assign z = ~a;
        end else begin : g_z_2
            // Preprocess a for increment/decrement
            assign at = a ^ {WIDTH{inc_dec}};

            // Calculate prefix output propagate signal
            AU_prefix_and #(
                .WIDTH(WIDTH),
                .ARCH (ARCH)
            ) u_AU_prefix_and (
                .pi(at),
                .po(po)
            );

            // Calculate result bits
            assign z = a ^ {po[WIDTH - 2 : 0], 1'b1};
        end
    endgenerate


endmodule
